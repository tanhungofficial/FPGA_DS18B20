library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity LCD_KHOI_TAO_HIEN_THI_FULL is
    Port (  LCD_DATA : out  STD_LOGIC_VECTOR (7 downto 0);
            LCD_RS, LCD_E : out  STD_LOGIC;
            LCD_CK, LCD_RST : in  STD_LOGIC;
			   H1_8:  in STD_LOGIC_VECTOR(7 DOWNTO 0);
				H1_9:  in STD_LOGIC_VECTOR(7 DOWNTO 0);
				H1_11: in STD_LOGIC_VECTOR(7 DOWNTO 0);	
				H1_12: in STD_LOGIC_VECTOR(7 DOWNTO 0);
				H1_14: in STD_LOGIC_VECTOR(7 DOWNTO 0);
				H1_15: in STD_LOGIC_VECTOR(7 DOWNTO 0);
				H2_11: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
				H2_12: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
				H2_13: IN STD_LOGIC_VECTOR(7 DOWNTO 0));
end LCD_KHOI_TAO_HIEN_THI_FULL;

architecture Behavioral of LCD_KHOI_TAO_HIEN_THI_FULL is
	-- KHAI BAO CAC BIEN 
TYPE LCD_MACHINE IS(
							LCD_INIT, 
							LCD_ADDR_L1,
							LCD_ADDR_L2,
							LCD_DATA_L1,
							LCD_DATA_L2,
							LCD_STOP	
							
							);
SIGNAL LCD_STATE: LCD_MACHINE:= LCD_INIT;
SIGNAL LCD_HANG_1,LCD_HANG_2: STD_LOGIC_VECTOR(127 DOWNTO 0);
TYPE LCD_CMD_TB IS ARRAY(INTEGER RANGE 0 TO 5) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
CONSTANT LCD_CMD : LCD_CMD_TB:= (
			0 =>  	X"00",
			1 =>  	X"3C", -- FUNCTION SET
			2 => 		X"0C", -- CONTROL DISPLAY
			3 => 		X"01", -- CLEAR
			4 => 		X"02", -- RETURN HOME
			5 => 		X"06"  -- ENTRY MODE SET
			);

TYPE LCD_DIS_L1 IS ARRAY(INTEGER RANGE 0 TO 15) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LCD_DIS1 : LCD_DIS_L1;

TYPE LCD_DIS_L2 IS ARRAY(INTEGER RANGE 0 TO 15) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL LCD_DIS2 : LCD_DIS_L2;

SIGNAL PTR : INTEGER RANGE 0 TO 15:=0;
SIGNAL SLX : INTEGER RANGE 0 TO 1000000 :=0;

BEGIN 
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= H1_8;
	LCD_HANG_1(79 DOWNTO 72)	<= H1_9;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(95 DOWNTO 88)	<= H1_11;
	LCD_HANG_1(103 DOWNTO 96)	<= H1_12;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(119 DOWNTO 112)	<= H1_14;
	LCD_HANG_1(127 DOWNTO 120)	<= H1_15;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(95 DOWNTO 88)	<= H2_11;
	LCD_HANG_2(103 DOWNTO 96)	<= H2_12;
	LCD_HANG_2(111 DOWNTO 104)	<= H2_13;
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('''),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	
	PROCESS(LCD_HANG_1,LCD_HANG_2)
	BEGIN
		FOR I IN 0 TO 15
		LOOP
			LCD_DIS1(I)<= LCD_HANG_1((I*8+7)DOWNTO I*8);
			LCD_DIS2(I)<= LCD_HANG_2((I*8+7)DOWNTO I*8);
		END LOOP;
	END PROCESS;
	
	PROCESS(LCD_CK,SLX,LCD_RST)
	BEGIN
		IF LCD_RST='1' THEN LCD_STATE					<= LCD_INIT;
								  SLX					<= 0;
								  PTR					<= 0;
								  
								 
		ELSIF	FALLING_EDGE(LCD_CK) THEN

			CASE LCD_STATE IS
				WHEN LCD_INIT => 		LCD_RS<='0';	
										SLX <= SLX + 1; 
					IF SLX = 164000 THEN	SLX <= 0;
						IF(PTR = 5 ) THEN   LCD_STATE <= LCD_ADDR_L1;
						ELSE 				PTR <= PTR + 1;
						END IF;
					ELSIF (SLX = 30) THEN LCD_E 	<= '0';
					ELSIF (SLX = 10) THEN LCD_E 	<= '1';
					ELSE		          LCD_DATA	<= LCD_CMD(PTR);					     	
					END IF;
				
				WHEN LCD_ADDR_L1 => 		LCD_RS<='0';
											SLX <= SLX + 1;
					IF SLX = 5000 THEN	SLX <= 0;
										LCD_STATE <= LCD_DATA_L1;
										PTR <= 0;
				
					ELSIF (SLX = 30) THEN LCD_E <= '0';
					ELSIF (SLX = 10) THEN LCD_E <= '1';
					ELSE
							LCD_DATA <=X"80";
					END IF;
												
				WHEN LCD_DATA_L1 => 		LCD_RS<='1';
											SLX <= SLX + 1;
					IF SLX = 5000 THEN		SLX <= 0;
						IF (PTR = 15) THEN 	LCD_STATE <= LCD_ADDR_L2;
						ELSE					  PTR <= PTR + 1;
						END IF;
					ELSIF (SLX = 30) THEN LCD_E <= '0';
					ELSIF (SLX = 10) THEN LCD_E <= '1';
					ELSE
							LCD_DATA <= LCD_DIS1(PTR);
					END IF;
				
				WHEN LCD_ADDR_L2 => 		LCD_RS<='0';
												SLX <= SLX + 1;
												IF SLX = 5000 THEN	SLX <= 0;
																					LCD_STATE <= LCD_DATA_L2;
																					PTR <= 0;
											
												ELSIF (SLX = 30) THEN LCD_E <= '0';
												ELSIF (SLX = 10) THEN LCD_E <= '1';
												ELSE
														LCD_DATA <=X"C0";
												END IF;
				WHEN LCD_DATA_L2 => 		LCD_RS<='1';
												SLX <= SLX + 1;
												IF SLX = 5000 THEN	SLX <= 0;
													IF (PTR = 15) THEN 	LCD_STATE <= LCD_STOP;
													ELSE									PTR <= PTR + 1;
													END IF;
												ELSIF (SLX = 30) THEN LCD_E <= '0';
												ELSIF (SLX = 10) THEN LCD_E <= '1';
												ELSE
														LCD_DATA <=  LCD_DIS2(PTR);
												END IF;
											  
				WHEN LCD_STOP	=> SLX <= SLX + 1;
										IF SLX = 1000000 THEN 	SLX <= 0;
																				LCD_STATE <= LCD_ADDR_L1;
										END IF;
				
				
			END CASE;
		END IF;						  
	END PROCESS;

end Behavioral;