library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;


entity LCD_KHOI_TAO_HIEN_THI_CGRAM_FULL is
PORT(	LCD_DB: 	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		LCD_RS,LCD_E: OUT STD_LOGIC;
		LCD_CK,LCD_RST: IN STD_LOGIC;
		H1_8:  in STD_LOGIC_VECTOR(7 DOWNTO 0);
		H1_9:  in STD_LOGIC_VECTOR(7 DOWNTO 0);
		H1_11: in STD_LOGIC_VECTOR(7 DOWNTO 0);	
		H1_12: in STD_LOGIC_VECTOR(7 DOWNTO 0);
		H1_14: in STD_LOGIC_VECTOR(7 DOWNTO 0);
		H1_15: in STD_LOGIC_VECTOR(7 DOWNTO 0);
		H2_11: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		H2_12: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		H2_13: IN STD_LOGIC_VECTOR(7 DOWNTO 0));
);
end LCD_KHOI_TAO_HIEN_THI_CGRAM_FULL;

architecture Behavioral of LCD_KHOI_TAO_HIEN_THI_CGRAM_FULL is
TYPE LCD_MACHINE IS(
							LCD_INITIAL,
							LCD_CGRAM_ADDRESS,
							LCD_CGRAM_DATA,
							LCD_ADDRESS_L1,
							LCD_DATA_L1,
							LCD_ADDRESS_L2,
							LCD_DATA_L2,
							LCD_STOP
);
SIGNAL LCD_HANG_1,LCD_HANG_2: STD_LOGIC_VECTOR(127 DOWNTO 0);
SIGNAL LCD_STATE: LCD_MACHINE:=LCD_INITIAL;
TYPE LCD_CMD_TABLE IS ARRAY (INTEGER RANGE 0 TO 5) OF STD_LOGIC_VECTOR(8 DOWNTO 0);
CONSTANT LCD_CMD: LCD_CMD_TABLE:=(0=> '0'&X"00",
                                  1=> '0'&X"3C",--FUNCTION SET
											 2=> '0'&X"0C",--DISLAY CONTROL
											 3=> '0'&X"01",--CLEAR
											 4=> '0'&X"02",--RETURN HOME
											 5=> '0'&X"06");--ENTRY MODE SET
SIGNAL LCD_CMD_PTR: INTEGER RANGE 0 TO 15:=0;

TYPE LCD_CGRAM_TABLE IS ARRAY (INTEGER RANGE 0 TO 63) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
CONSTANT LCD_CGRAM: LCD_CGRAM_TABLE:= (
	X"07", X"0F", X"1F", X"1F", X"1F", X"1F", X"1F", X"1F",---F-0
	X"1F", X"1F", X"1F", X"00", X"00", X"00", X"00", X"00",---A-1
	X"1C", X"1E", X"1F", X"1F", X"1F", X"1F", X"1F", X"1F",---B-2
	X"00", X"00", X"00", X"00", X"00", X"1F", X"1F", X"1F",---D-3
	X"1F", X"1F", X"1F", X"1F", X"1F", X"1F", X"1E", X"1C",---C-4
	X"1F", X"1F", X"1F", X"1F", X"1F", X"1F", X"0F", X"07",---E-5
	X"1F", X"1F", X"1F", X"00", X"00", X"00", X"1F", X"1F",---G+D-6
	X"1F", X"1F", X"1F", X"1F", X"1F", X"1F", X"1F", X"1F"---I-7
); 


SIGNAL LCD_CGRAM_PTR: INTEGER RANGE 0 TO LCD_CGRAM'HIGH:=0;

TYPE 	LCD_DIS_L1 IS ARRAY (INTEGER RANGE 0 TO 15) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL 	LCD_DIS1:LCD_DIS_L1;
TYPE 	LCD_DIS_L2 IS ARRAY (INTEGER RANGE 0 TO 15) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL 	LCD_DIS2:LCD_DIS_L2;
SIGNAL 	LCD_DIS_PTR: INTEGER RANGE 0 TO 15:=0;
SIGNAL 	LCD_DELAY: INTEGER RANGE 0 TO 1000000:=0;
SIGNAL 	LCD_RS_DB: STD_LOGIC_VECTOR(8 DOWNTO 0):='0'&X"00";
SIGNAL 	LCD_ENABLE: STD_LOGIC:='0';
begin
//	GAN DU LIEU

	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= H1_8;
	LCD_HANG_1(79 DOWNTO 72)	<= H1_9;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(95 DOWNTO 88)	<= H1_11;
	LCD_HANG_1(103 DOWNTO 96)	<= H1_12;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(119 DOWNTO 112)	<= H1_14;
	LCD_HANG_1(127 DOWNTO 120)	<= H1_15;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(95 DOWNTO 88)	<= H2_11;
	LCD_HANG_2(103 DOWNTO 96)	<= H2_12;
	LCD_HANG_2(111 DOWNTO 104)	<= H2_13;
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('''),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	
	
  PROCESS(LCD_HANG_1,LCD_HANG_2)
  BEGIN
    FOR I IN 0 TO 15
	 LOOP
	     LCD_DIS1(I) <=LCD_HANG_1((I*8+7) DOWNTO I*8);
        LCD_DIS2(I) <=LCD_HANG_2((I*8+7) DOWNTO I*8);
	 END LOOP;
  END PROCESS;
  
  PROCESS(LCD_CK,LCD_DELAY,LCD_RST)
  BEGIN
  IF LCD_RST='1' THEN LCD_STATE<=LCD_INITIAL;
                      LCD_DELAY<=0;
							 LCD_CMD_PTR<=0;
							 LCD_DIS_PTR<=0;
							 LCD_CGRAM_PTR <= 0;
	ELSIF FALLING_EDGE(LCD_CK) THEN
	   CASE LCD_STATE IS
		  WHEN LCD_INITIAL=>  LCD_DELAY<=LCD_DELAY+1;
		                      IF LCD_DELAY = 164000 THEN LCD_DELAY<=0;
									    IF (LCD_CMD_PTR= LCD_CMD'HIGH) THEN 
										                                       LCD_STATE<=LCD_CGRAM_ADDRESS;
											ELSE	
                                    											LCD_CMD_PTR<=LCD_CMD_PTR+1;
											END IF;
									ELSIF(LCD_DELAY=30) THEN LCD_ENABLE<='0';
									ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									ELSE                     LCD_RS_DB<=LCD_CMD(LCD_CMD_PTR);
									END IF;
			WHEN LCD_CGRAM_ADDRESS => LCD_DELAY<=LCD_DELAY+1;
		                       IF LCD_DELAY=5000 THEN LCD_DELAY<=0;
									                         LCD_STATE<=LCD_CGRAM_DATA;
																	 LCD_DIS_PTR<=0;
									  ELSIF (LCD_DELAY=30)THEN LCD_ENABLE<='0';
								     ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									  ELSE                     LCD_RS_DB<='0'&X"40";
									  END IF;
			WHEN LCD_CGRAM_DATA=>    LCD_DELAY<=LCD_DELAY+1;
		                      IF LCD_DELAY=5000 THEN LCD_DELAY<=0;
									    IF (LCD_CGRAM_PTR= LCD_CGRAM'HIGH) THEN 
										                                       LCD_STATE<=LCD_ADDRESS_L1;
											ELSE	
                                    											LCD_CGRAM_PTR<=LCD_CGRAM_PTR+1;
											END IF;
									ELSIF(LCD_DELAY=30) THEN LCD_ENABLE<='0';
									ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									ELSE                     LCD_RS_DB<='1'& LCD_CGRAM(LCD_CGRAM_PTR);
									END IF;				
		 WHEN LCD_ADDRESS_L1=> LCD_DELAY<=LCD_DELAY+1;
		                       IF LCD_DELAY=5000 THEN 	LCD_DELAY<=0;
									                    LCD_STATE<=LCD_DATA_L1;
														LCD_DIS_PTR<=0;
									  ELSIF (LCD_DELAY=30)THEN LCD_ENABLE<='0';
								     ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									  ELSE                     LCD_RS_DB<='0'&X"80";
									  END IF;
		WHEN LCD_DATA_L1=>    LCD_DELAY<=LCD_DELAY+1;
		                      IF LCD_DELAY=5000 THEN LCD_DELAY<=0;
									    IF (LCD_DIS_PTR=15) THEN LCD_STATE<=LCD_ADDRESS_L2;
										 ELSE                     LCD_DIS_PTR<=LCD_DIS_PTR+1;
										 END IF;
									ELSIF(LCD_DELAY=30) THEN LCD_ENABLE<='0';
									ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									ELSE                     LCD_RS_DB<='1'& LCD_DIS1(LCD_DIS_PTR);
									END IF;
		WHEN LCD_ADDRESS_L2=> LCD_DELAY<=LCD_DELAY+1;
		                       IF LCD_DELAY=5000 THEN LCD_DELAY<=0;
																	LCD_STATE<=LCD_DATA_L2;
																	LCD_DIS_PTR<=0;
									  ELSIF (LCD_DELAY=30)THEN 	LCD_ENABLE<='0';
								     ELSIF(LCD_DELAY=5)  THEN 	LCD_ENABLE<='1';
									  ELSE                     	LCD_RS_DB<='0'&X"C0";
									  END IF;
		WHEN LCD_DATA_L2=>    LCD_DELAY<=LCD_DELAY+1;
		                      IF LCD_DELAY=5000 THEN LCD_DELAY<=0;
									    IF (LCD_DIS_PTR=15) THEN LCD_STATE<=LCD_STOP;
										 ELSE                    LCD_DIS_PTR<=LCD_DIS_PTR+1;
										 END IF;
									ELSIF(LCD_DELAY=30) THEN LCD_ENABLE<='0';
									ELSIF(LCD_DELAY=5)  THEN LCD_ENABLE<='1';
									ELSE                     LCD_RS_DB<='1'& LCD_DIS2(LCD_DIS_PTR);
									END IF;
	   WHEN LCD_STOP=>    LCD_DELAY<=LCD_DELAY+1;
		                   IF LCD_DELAY=1000000 THEN 		LCD_DELAY<=0;
															LCD_STATE<=LCD_ADDRESS_L1;
								END IF;
		END CASE;
	END IF;
  END PROCESS;
  LCD_DB<=LCD_RS_DB( 7 DOWNTO 0);
  LCD_RS<=LCD_RS_DB(8);
  LCD_E<=LCD_ENABLE;
end Behavioral;

